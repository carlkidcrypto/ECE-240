`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:14:41 03/05/2019 
// Design Name: 
// Module Name:    comparator_2b 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module comparator_2b(A, B, G, L, E);
    input [2:0] A;
    input [2:0] B;
    output [2:0] G;
    output [2:0] L;
    output [2:0] E;


endmodule
