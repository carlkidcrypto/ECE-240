`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:35:42 03/25/2019 
// Design Name: 
// Module Name:    Crazy_Counter_up1_dwn2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Crazy_Counter_up1_dwn2(CLK, RST, cnt, cnt_dir, load_enb);
    input CLK;
    input RST;
    output [3:0] cnt;
    input cnt_dir;
    input load_enb;


endmodule
